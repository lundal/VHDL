library IEEE;
use IEEE.STD_LOGIC_1164.ALL;

entity memory_stage is
end memory_stage;

architecture Behavioral of memory_stage is

begin


end Behavioral;

