library IEEE;
use IEEE.STD_LOGIC_1164.ALL;

entity write_back_stage is
end write_back_stage;

architecture Behavioral of write_back_stage is

begin


end Behavioral;

